
function [255:0] bram_ini_table;
input integer index;//Mode type 
input integer val_; //Port A index, Port B Index, Number of Items in Loop, Port A Start, Port B Start, reserved 
case (index)
   0: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
   1: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
   2: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
   3: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
   4: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
   5: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
   6: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
   7: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
   8: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
   9: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  10: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  11: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  12: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  13: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  14: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  15: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  16: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  17: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  18: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  19: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  20: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  21: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  22: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  23: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  24: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  25: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  26: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  27: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  28: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  29: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  30: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  31: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  32: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  33: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  34: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  35: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  36: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  37: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  38: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  39: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  40: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  41: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  42: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  43: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  44: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  45: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  46: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  47: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  48: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  49: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  50: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
  51: bram_ini_table=
(val_== 0)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 1)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 2)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 3)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 4)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 5)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 6)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 7)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 8)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_== 9)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==10)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==11)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==12)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==13)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==14)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==15)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==16)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==17)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==18)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==19)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==20)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==21)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==22)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==23)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==24)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==25)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==26)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==27)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==28)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==29)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==30)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==31)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==32)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==33)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==34)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==35)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==36)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==37)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==38)?256'h0000000000000000000000000000000000000000000000000000000000000000:
(val_==39)?256'h0000000000000000000000000000000000000000000000000000000000000000:
0;
   endcase
endfunction  
